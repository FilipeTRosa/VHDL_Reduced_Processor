library ieee;                 
use ieee.std_logic_1164.all;  
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

entity decod8x256 is 
	port(
		endereco	: in std_logic_vector(7 downto 0);
		saida		: out integer
	);
end entity;
architecture behavior of decod8x256 is 
begin

	saida <= 0   when endereco = "00000000" else
             1   when endereco = "00000001" else
             2   when endereco = "00000010" else
             3   when endereco = "00000011" else
             4   when endereco = "00000100" else
             5   when endereco = "00000101" else
             6   when endereco = "00000110" else
             7   when endereco = "00000111" else
             8   when endereco = "00001000" else
             9   when endereco = "00001001" else
             10  when endereco = "00001010" else
             11  when endereco = "00001011" else
             12  when endereco = "00001100" else
             13  when endereco = "00001101" else
             14  when endereco = "00001110" else
             15  when endereco = "00001111" else
             16  when endereco = "00010000" else
             17  when endereco = "00010001" else
             18  when endereco = "00010010" else
             19  when endereco = "00010011" else
             20  when endereco = "00010100" else
             21  when endereco = "00010101" else
             22  when endereco = "00010110" else
             23  when endereco = "00010111" else
             24  when endereco = "00011000" else
             25  when endereco = "00011001" else
             26  when endereco = "00011010" else
             27  when endereco = "00011011" else
             28  when endereco = "00011100" else
             29  when endereco = "00011101" else
             30  when endereco = "00011110" else
             31  when endereco = "00011111" else
             32  when endereco = "00100000" else
             33  when endereco = "00100001" else
             34  when endereco = "00100010" else
             35  when endereco = "00100011" else
             36  when endereco = "00100100" else
             37  when endereco = "00100101" else
             38  when endereco = "00100110" else
             39  when endereco = "00100111" else
             40  when endereco = "00101000" else
             41  when endereco = "00101001" else
             42  when endereco = "00101010" else
             43  when endereco = "00101011" else
             44  when endereco = "00101100" else
             45  when endereco = "00101101" else
             46  when endereco = "00101110" else
             47  when endereco = "00101111" else
             48  when endereco = "00110000" else
             49  when endereco = "00110001" else
             50  when endereco = "00110010" else
             51  when endereco = "00110011" else
             52  when endereco = "00110100" else
             53  when endereco = "00110101" else
             54  when endereco = "00110110" else
             55  when endereco = "00110111" else
             56  when endereco = "00111000" else
             57  when endereco = "00111001" else
             58  when endereco = "00111010" else
             59  when endereco = "00111011" else
             60  when endereco = "00111100" else
             61  when endereco = "00111101" else
             62  when endereco = "00111110" else
             63  when endereco = "00111111" else
             64  when endereco = "01000000" else
             65  when endereco = "01000001" else
             66  when endereco = "01000010" else
             67  when endereco = "01000011" else
             68  when endereco = "01000100" else
             69  when endereco = "01000101" else
             70  when endereco = "01000110" else
             71  when endereco = "01000111" else
             72  when endereco = "01001000" else
             73  when endereco = "01001001" else
             74  when endereco = "01001010" else
             75  when endereco = "01001011" else
             76  when endereco = "01001100" else
             77  when endereco = "01001101" else
             78  when endereco = "01001110" else
             79  when endereco = "01001111" else
             80  when endereco = "01010000" else
             81  when endereco = "01010001" else
             82  when endereco = "01010010" else
             83  when endereco = "01010011" else
             84  when endereco = "01010100" else
             85  when endereco = "01010101" else
             86  when endereco = "01010110" else
             87  when endereco = "01010111" else
             88  when endereco = "01011000" else
             89  when endereco = "01011001" else
             90  when endereco = "01011010" else
             91  when endereco = "01011011" else
             92  when endereco = "01011100" else
             93  when endereco = "01011101" else
             94  when endereco = "01011110" else
             95  when endereco = "01011111" else
             96  when endereco = "01100000" else
             97  when endereco = "01100001" else
             98  when endereco = "01100010" else
             99  when endereco = "01100011" else
             100 when endereco = "01100100" else
             101 when endereco = "01100101" else
             102 when endereco = "01100110" else
             103 when endereco = "01100111" else
             104 when endereco = "01101000" else
             105 when endereco = "01101001" else
             106 when endereco = "01101010" else
             107 when endereco = "01101011" else
             108 when endereco = "01101100" else
             109 when endereco = "01101101" else
             110 when endereco = "01101110" else
             111 when endereco = "01101111" else
             112 when endereco = "01110000" else
             113 when endereco = "01110001" else
             114 when endereco = "01110010" else
             115 when endereco = "01110011" else
             116 when endereco = "01110100" else
             117 when endereco = "01110101" else
             118 when endereco = "01110110" else
             119 when endereco = "01110111" else
             120 when endereco = "01111000" else
             121 when endereco = "01111001" else
             122 when endereco = "01111010" else
             123 when endereco = "01111011" else
             124 when endereco = "01111100" else
             125 when endereco = "01111101" else
             126 when endereco = "01111110" else
             127 when endereco = "01111111" else
             128 when endereco = "10000000" else
             129 when endereco = "10000001" else
             130 when endereco = "10000010" else
             131 when endereco = "10000011" else
             132 when endereco = "10000100" else
             133 when endereco = "10000101" else
             134 when endereco = "10000110" else
             135 when endereco = "10000111" else
             136 when endereco = "10001000" else
             137 when endereco = "10001001" else
             138 when endereco = "10001010" else
             139 when endereco = "10001011" else
             140 when endereco = "10001100" else
             141 when endereco = "10001101" else
             142 when endereco = "10001110" else
             143 when endereco = "10001111" else
             144 when endereco = "10010000" else
             145 when endereco = "10010001" else
             146 when endereco = "10010010" else
             147 when endereco = "10010011" else
             148 when endereco = "10010100" else
             149 when endereco = "10010101" else
             150 when endereco = "10010110" else
             151 when endereco = "10010111" else
             152 when endereco = "10011000" else
             153 when endereco = "10011001" else
             154 when endereco = "10011010" else
             155 when endereco = "10011011" else
             156 when endereco = "10011100" else
             157 when endereco = "10011101" else
             158 when endereco = "10011110" else
             159 when endereco = "10011111" else
             160 when endereco = "10100000" else
             161 when endereco = "10100001" else
             162 when endereco = "10100010" else
             163 when endereco = "10100011" else
             164 when endereco = "10100100" else
             165 when endereco = "10100101" else
             166 when endereco = "10100110" else
             167 when endereco = "10100111" else
             168 when endereco = "10101000" else
             169 when endereco = "10101001" else
             170 when endereco = "10101010" else
             171 when endereco = "10101011" else
             172 when endereco = "10101100" else
             173 when endereco = "10101101" else
             174 when endereco = "10101110" else
             175 when endereco = "10101111" else
             176 when endereco = "10110000" else
             177 when endereco = "10110001" else
             178 when endereco = "10110010" else
             179 when endereco = "10110011" else
             180 when endereco = "10110100" else
             181 when endereco = "10110101" else
             182 when endereco = "10110110" else
             183 when endereco = "10110111" else
             184 when endereco = "10111000" else
             185 when endereco = "10111001" else
             186 when endereco = "10111010" else
             187 when endereco = "10111011" else
             188 when endereco = "10111100" else
             189 when endereco = "10111101" else
             190 when endereco = "10111110" else
             191 when endereco = "10111111" else
             192 when endereco = "11000000" else
             193 when endereco = "11000001" else
             194 when endereco = "11000010" else
             195 when endereco = "11000011" else
             196 when endereco = "11000100" else
             197 when endereco = "11000101" else
             198 when endereco = "11000110" else
             199 when endereco = "11000111" else
             200 when endereco = "11001000" else
             201 when endereco = "11001001" else
             202 when endereco = "11001010" else
             203 when endereco = "11001011" else
             204 when endereco = "11001100" else
             205 when endereco = "11001101" else
             206 when endereco = "11001110" else
             207 when endereco = "11001111" else
             208 when endereco = "11010000" else
             209 when endereco = "11010001" else
             210 when endereco = "11010010" else
             211 when endereco = "11010011" else
             212 when endereco = "11010100" else
             213 when endereco = "11010101" else
             214 when endereco = "11010110" else
             215 when endereco = "11010111" else
             216 when endereco = "11011000" else
             217 when endereco = "11011001" else
             218 when endereco = "11011010" else
             219 when endereco = "11011011" else
             220 when endereco = "11011100" else
             221 when endereco = "11011101" else
             222 when endereco = "11011110" else
             223 when endereco = "11011111" else
             224 when endereco = "11100000" else
             225 when endereco = "11100001" else
             226 when endereco = "11100010" else
             227 when endereco = "11100011" else
             228 when endereco = "11100100" else
             229 when endereco = "11100101" else
             230 when endereco = "11100110" else
             231 when endereco = "11100111" else
             232 when endereco = "11101000" else
             233 when endereco = "11101001" else
             234 when endereco = "11101010" else
             235 when endereco = "11101011" else
             236 when endereco = "11101100" else
             237 when endereco = "11101101" else
             238 when endereco = "11101110" else
             239 when endereco = "11101111" else
             240 when endereco = "11110000" else
             241 when endereco = "11110001" else
             242 when endereco = "11110010" else
             243 when endereco = "11110011" else
             244 when endereco = "11110100" else
             245 when endereco = "11110101" else
             246 when endereco = "11110110" else
             247 when endereco = "11110111" else
             248 when endereco = "11111000" else
             249 when endereco = "11111001" else
             250 when endereco = "11111010" else
             251 when endereco = "11111011" else
             252 when endereco = "11111100" else
             253 when endereco = "11111101" else
             254 when endereco = "11111110" else
             255 when endereco = "11111111";

end behavior;